`timescale 1ns / 1ps
//fdivider_10.v
module freq_divider_by_10 #(
    parameter DIVISOR = 10
)(
    input wire clk_in,
    input wire reset,
    output reg clk_out
);

endmodule
