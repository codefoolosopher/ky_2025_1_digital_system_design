
`timescale 1ns / 1ps

module shift_register_sipo #(
    parameter WIDTH = 8
)(
    input clk,
    input reset,
    input serial_in,
    output reg [7:0] parallel_out
);


endmodule
