`timescale 1ns / 1ps
module Testbench;

    reg clk;
    reg reset;
    reg write_enable;
    reg [7:0] write_data;
    wire [7:0] read_data;


endmodule
