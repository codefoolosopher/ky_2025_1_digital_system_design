`timescale 1ns / 1ps
module seq_detector_1010(input clk, rst_n, x, output reg z);
  parameter A = 4'h1;
  parameter B = 4'h2;
  parameter C = 4'h3;
  parameter D = 4'h4;
  parameter E = 4'h5; // extra state when compared with Mealy Machine
  
endmodule